magic
tech sky130A
magscale 1 2
timestamp 1740936470
<< locali >>
rect -82 -1742 110 -1478
rect 1072 -1742 1264 -1458
rect -130 -1756 1288 -1742
rect -130 -1934 312 -1756
rect 492 -1934 1288 -1756
<< viali >>
rect 312 -1936 492 -1756
<< metal1 >>
rect 178 740 242 2246
rect 690 2156 1148 2348
rect 240 676 242 740
rect 178 -1566 242 676
rect 306 -1756 498 1960
rect 956 1558 1148 2156
rect 684 1366 1148 1558
rect 742 740 806 746
rect 742 670 806 676
rect 956 -58 1148 1366
rect 688 -250 1148 -58
rect 688 -618 880 -376
rect 956 -1074 1148 -250
rect 688 -1266 1148 -1074
rect 306 -1936 312 -1756
rect 492 -1936 498 -1756
rect 306 -1948 498 -1936
<< via1 >>
rect 176 676 240 740
rect 764 676 868 740
<< metal2 >>
rect -145 740 789 741
rect -146 676 176 740
rect 240 676 764 740
rect 868 676 874 740
rect -145 675 789 676
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ~/pro/aicex/ip/jnw_ex_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 16 0 1 24
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1734044400
transform 1 0 14 0 1 834
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1734044400
transform 1 0 16 0 1 -794
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1734044400
transform 1 0 18 0 1 1656
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_5
timestamp 1734044400
transform 1 0 16 0 1 -1610
box -184 -128 1336 928
<< labels >>
flabel metal2 -146 676 -82 740 0 FreeSans 8 0 0 0 IBPS_5U
flabel metal2 -144 676 -80 740 0 FreeSans 1600 0 0 0 IBPS_5U
flabel metal1 956 676 1148 868 0 FreeSans 1600 0 0 0 IBNS_20U
flabel viali 312 -1936 492 -1756 0 FreeSans 1600 0 0 0 VSS
<< end >>
